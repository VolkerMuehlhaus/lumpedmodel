* EQUIVALENT CIRCUIT FOR VECTOR FITTED S-MATRIX
* Created using scikit-rf vectorFitting.py
*
.SUBCKT s_equivalent p1 p2
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 0.0042024138934587925
Fd1_1 0 s1 V1 0.21012069467293965
Gr1_re_1_1 0 s1 x1_re_a1 0 -79045098281.26822
Gr1_im_1_1 0 s1 x1_im_a1 0 -55444207716.82171
Gr2_1_1 0 s1 x2_a1 0 -10024001.170605147
Gr3_1_1 0 s1 x3_a1 0 -10345375682.877348
Gr4_1_1 0 s1 x4_a1 0 462193161579.34717
Gr5_1_1 0 s1 x5_a1 0 -278458975143.8581
Gd1_2 0 s1 p2 0 0.007706882576195599
Fd1_2 0 s1 V2 0.38534412880978
Gr1_re_1_2 0 s1 x1_re_a2 0 -27235147402.452938
Gr1_im_1_2 0 s1 x1_im_a2 0 4326911607.167198
Gr2_1_2 0 s1 x2_a2 0 40912942.50726339
Gr3_1_2 0 s1 x3_a2 0 10527646259.764256
Gr4_1_2 0 s1 x4_a2 0 -387896015833.9557
Gr5_1_2 0 s1 x5_a2 0 268583538097.7818
*
* State networks driven by port 1
Cx1_re_a1 x1_re_a1 0 1.0
Gx1_re_a1 0 x1_re_a1 p1 0 0.1414213562373095
Fx1_re_a1 0 x1_re_a1 V1 7.0710678118654755
Rp1_re_re_a1 0 x1_re_a1 3.3680980971317083e-12
Gp1_re_im_a1 0 x1_re_a1 x1_im_a1 0 926824465249.058
Cx1_im_a1 x1_im_a1 0 1.0
Gp1_im_re_a1 0 x1_im_a1 x1_re_a1 0 -926824465249.058
Rp1_im_im_a1 0 x1_im_a1 3.3680980971317083e-12
Cx2_a1 x2_a1 0 1.0
Gx2_a1 0 x2_a1 p1 0 0.07071067811865475
Fx2_a1 0 x2_a1 V1 3.5355339059327378
Rp2_a1 0 x2_a1 5.884474762399651e-11
Cx3_a1 x3_a1 0 1.0
Gx3_a1 0 x3_a1 p1 0 0.07071067811865475
Fx3_a1 0 x3_a1 V1 3.5355339059327378
Rp3_a1 0 x3_a1 5.772531776779665e-12
Cx4_a1 x4_a1 0 1.0
Gx4_a1 0 x4_a1 p1 0 0.07071067811865475
Fx4_a1 0 x4_a1 V1 3.5355339059327378
Rp4_a1 0 x4_a1 1.3813640211512772e-12
Cx5_a1 x5_a1 0 1.0
Gx5_a1 0 x5_a1 p1 0 0.07071067811865475
Fx5_a1 0 x5_a1 V1 3.5355339059327378
Rp5_a1 0 x5_a1 2.486019786956729e-12
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 0.007706882591895254
Fd2_1 0 s2 V1 0.3853441295947627
Gr1_re_2_1 0 s2 x1_re_a1 0 -27235147458.442665
Gr1_im_2_1 0 s2 x1_im_a1 0 4326911552.570392
Gr2_2_1 0 s2 x2_a1 0 40912945.409499735
Gr3_2_1 0 s2 x3_a1 0 10527646229.574852
Gr4_2_1 0 s2 x4_a1 0 -387896016337.9314
Gr5_2_1 0 s2 x5_a1 0 268583538316.9227
Gd2_2 0 s2 p2 0 0.0034053893291790347
Fd2_2 0 s2 V2 0.17026946645895175
Gr1_re_2_2 0 s2 x1_re_a2 0 -69230643064.64342
Gr1_im_2_2 0 s2 x1_im_a2 0 -54811433523.57486
Gr2_2_2 0 s2 x2_a2 0 -9674637.488665758
Gr3_2_2 0 s2 x3_a2 0 -10261904844.476898
Gr4_2_2 0 s2 x4_a2 0 461564904098.4481
Gr5_2_2 0 s2 x5_a2 0 -275760684961.0225
*
* State networks driven by port 2
Cx1_re_a2 x1_re_a2 0 1.0
Gx1_re_a2 0 x1_re_a2 p2 0 0.1414213562373095
Fx1_re_a2 0 x1_re_a2 V2 7.0710678118654755
Rp1_re_re_a2 0 x1_re_a2 3.3680980971317083e-12
Gp1_re_im_a2 0 x1_re_a2 x1_im_a2 0 926824465249.058
Cx1_im_a2 x1_im_a2 0 1.0
Gp1_im_re_a2 0 x1_im_a2 x1_re_a2 0 -926824465249.058
Rp1_im_im_a2 0 x1_im_a2 3.3680980971317083e-12
Cx2_a2 x2_a2 0 1.0
Gx2_a2 0 x2_a2 p2 0 0.07071067811865475
Fx2_a2 0 x2_a2 V2 3.5355339059327378
Rp2_a2 0 x2_a2 5.884474762399651e-11
Cx3_a2 x3_a2 0 1.0
Gx3_a2 0 x3_a2 p2 0 0.07071067811865475
Fx3_a2 0 x3_a2 V2 3.5355339059327378
Rp3_a2 0 x3_a2 5.772531776779665e-12
Cx4_a2 x4_a2 0 1.0
Gx4_a2 0 x4_a2 p2 0 0.07071067811865475
Fx4_a2 0 x4_a2 V2 3.5355339059327378
Rp4_a2 0 x4_a2 1.3813640211512772e-12
Cx5_a2 x5_a2 0 1.0
Gx5_a2 0 x5_a2 p2 0 0.07071067811865475
Fx5_a2 0 x5_a2 V2 3.5355339059327378
Rp5_a2 0 x5_a2 2.486019786956729e-12
.ENDS s_equivalent
